* start of a spice file
.model blah
.start
R3 vcc 5V 1.05368521445554K
R1 vcc intb 10.0mEG
R2 intb 0 100.0m RESMOD
CoUT out 5V 10u
Cin intb in 10000.0n
C2 intb in 4.7u
C3 intb in 1000n
M1 intb in 5V 0 pmos
pfet1 intb 0 5V inta in modelname
x1234 out inta in intb 0 modelname

.commands
.end
 
.

