* start of a spice file
.model blah
.start
R3 vcc 5V 1.0K
R1 vcc intb 10.0mEG
R2 intb 0 100.0m RESMOD
Cout out 5V 10u
Cin intb in 10000.0n
C2 intb in 4.7u
C3 intb in 1000n
M1 intb in 5V 0 pmos
.commands
.end
 
.

